library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std;


entity result is
        PORT (ledIN : IN BIT_VECTOR (2 downto 0);
               r : IN BIT_VECTOR (1 downto 0);
               buttons : IN BIT_VECTOR (2 downto 0);
               result : OUT BIT_VECTOR (2 downto 0));
end result;


architecture behavior of result is
begin
  process (ledIN,r,buttons)
  begin
	  if (buttons = "100") then
		result <= buttons;
	  elsif (buttons = "010") then
		result <= buttons;
	  elsif (buttons = "001") then
		result <= buttons;
	  elsif (r = "00") then
		result <= ledIN;
	  elsif (r = "01") then
		result <= (ledIN ror 1);
	  elsif (r = "10") then
		result <= (ledIN rol 1);
	  else
		result <= ledIN;
	  end if;
  end process;
  
end behavior;